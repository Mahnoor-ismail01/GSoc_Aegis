```
import uvm_pkg::*;
`include "adder_add_operation_packet.sv"

class adder_reset_test_seq extends uvm_sequence;
  `uvm_object_utils(adder_reset_test_seq)

  // Reference to the transaction packet
  rand adder_add_operation_packet pkt;

  // Constructor
  function new(string name = "adder_reset_test_seq");
    super.new(name);
  endfunction

  // Body task to generate and randomize transactions
  virtual task body();
    repeat (5) begin
      `uvm_info("SEQUENCE", $sformatf("Starting iteration %0d for %s", this.get_sequence_id(), "reset_test"), UVM_LOW)
      pkt = adder_add_operation_packet::type_id::create("pkt");
      if (!pkt.randomize() with {
        
        rstn == 0;
        
      }) begin
        `uvm_error("RANDOMIZE", "Randomization failed")
      end

      // Apply delay
      #50;

      // Start item and finish item
      start_item(pkt);
      finish_item(pkt);

      // Check expected output (basic comparison)
      if (pkt.rstn) begin
        if (pkt.sum != (pkt.a + pkt.b)[7:0] || pkt.carry != (pkt.a + pkt.b)[8]) begin
          `uvm_error("CHECK", $sformatf("Mismatch: sum=%0h, carry=%0b, expected sum=%0h, carry=%0b", pkt.sum, pkt.carry, (pkt.a + pkt.b)[7:0], (pkt.a + pkt.b)[8]))
        end
      
        if (pkt.sum != 0) begin
          `uvm_error("CHECK", $sformatf("Expected sum=%s, got %s", 0, pkt.sum))
        end
      
        if (pkt.carry != 0) begin
          `uvm_error("CHECK", $sformatf("Expected carry=%s, got %s", 0, pkt.carry))
        end
      
      end else begin
        if (pkt.sum != 0 || pkt.carry != 0) begin
          `uvm_error("CHECK", "Reset active but sum or carry not zero")
        end
      end
    end
  endtask
endclass
```