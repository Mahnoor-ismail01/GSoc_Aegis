
class corner_case_max_sequence extends uvm_sequence #(adder_transaction);
  `uvm_object_utils(corner_case_max_sequence)
  
  function new(string name = "corner_case_max_sequence");
    super.new(name);
  endfunction
  
  task body();
    adder_transaction tx;
    
    tx = adder_transaction::type_id::create("tx");
    start_item(tx);
    finish_item(tx);
    
  endtask
endclass